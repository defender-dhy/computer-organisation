`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:04:57 09/02/2020 
// Design Name: 
// Module Name:    add 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module add(input[7:0]a ,input[4:7]b,input[7:0]c,output[7:0] result);
wire w1, w2;
reg r1, r2;

assign r1=w1;
assign r1=r1+1;
endmodule

module AndGate(input[7:0] a,input[7:0] b,input[7:0] c,output[7:0] result);

    assign C=temp?B:A;

endmodule